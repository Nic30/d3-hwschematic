module constPortDriver(output out);
  assign out = 1;
endmodule

