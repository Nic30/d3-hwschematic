module subModuleBlackbox(output out);
  subSubModuleBlackbox b(out);
endmodule

