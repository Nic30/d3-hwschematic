module constAdder(input [8-1:0] in, output [8-1:0] out);
  assign out = in + 8'B 10101101;
endmodule
