module split1(input [8-1:0] in, output [4-1:0] out);
  assign out = in[5-1:1];
endmodule
