module subModuleBlackbox2(output out);
  subSubModuleBlackbox b(out);
endmodule

