module wireModule(input [8-1:0] in, output [8-1:0] out);
  assign out = in;
endmodule
